magic
tech scmos
timestamp 1427389379
<< pwell >>
rect -39 -45 23 -2
<< nwell >>
rect -39 2 23 65
<< polysilicon >>
rect -4 62 -2 64
rect 6 62 8 64
rect -24 25 -22 28
rect -4 25 -2 42
rect 6 39 8 42
rect 6 25 8 35
rect -24 -5 -22 5
rect -4 -5 -2 5
rect 6 -5 8 5
rect -24 -18 -22 -15
rect -4 -25 -2 -15
rect -4 -32 -2 -29
rect 6 -32 8 -15
rect -4 -44 -2 -42
rect 6 -44 8 -42
<< ndiffusion >>
rect -26 -15 -24 -5
rect -22 -15 -20 -5
rect -6 -15 -4 -5
rect -2 -15 0 -5
rect 4 -15 6 -5
rect 8 -15 10 -5
rect -6 -42 -4 -32
rect -2 -42 0 -32
rect 4 -42 6 -32
rect 8 -42 10 -32
<< pdiffusion >>
rect -6 42 -4 62
rect -2 42 0 62
rect 4 42 6 62
rect 8 42 10 62
rect -26 5 -24 25
rect -22 5 -20 25
rect -6 5 -4 25
rect -2 5 0 25
rect 4 5 6 25
rect 8 5 10 25
<< metal1 >>
rect -51 65 -32 69
rect -28 65 33 69
rect -25 64 -21 65
rect 0 62 4 65
rect -51 42 -15 46
rect -11 42 -10 62
rect 14 42 15 62
rect 22 42 33 46
rect 22 39 26 42
rect -39 35 2 39
rect 9 35 26 39
rect -39 2 -35 35
rect -2 32 2 35
rect -21 28 -6 32
rect -2 28 14 32
rect -32 25 -28 28
rect -10 25 -6 28
rect 10 25 14 28
rect -32 5 -30 25
rect -20 2 -16 5
rect -39 -2 -16 2
rect -20 -5 -16 -2
rect 0 2 4 5
rect 0 -2 23 2
rect 0 -5 4 -2
rect -31 -15 -30 -5
rect -16 -15 -10 -5
rect 10 -18 14 -15
rect -39 -22 -25 -18
rect -21 -22 14 -18
rect -1 -29 15 -25
rect -11 -42 -10 -32
rect 14 -42 15 -32
rect -26 -45 -22 -44
rect 0 -45 4 -42
rect -51 -49 -35 -45
rect -31 -49 33 -45
<< metal2 >>
rect -43 -18 -39 75
rect -32 32 -28 65
rect -35 -45 -31 -15
rect -15 -32 -11 42
rect 15 -25 19 42
rect 15 -32 19 -29
rect 23 -49 27 -2
<< ntransistor >>
rect -24 -15 -22 -5
rect -4 -15 -2 -5
rect 6 -15 8 -5
rect -4 -42 -2 -32
rect 6 -42 8 -32
<< ptransistor >>
rect -4 42 -2 62
rect 6 42 8 62
rect -24 5 -22 25
rect -4 5 -2 25
rect 6 5 8 25
<< polycontact >>
rect -25 28 -21 32
rect 5 35 9 39
rect -25 -22 -21 -18
rect -5 -29 -1 -25
<< ndcontact >>
rect -30 -15 -26 -5
rect -20 -15 -16 -5
rect -10 -15 -6 -5
rect 0 -15 4 -5
rect 10 -15 14 -5
rect -10 -42 -6 -32
rect 0 -42 4 -32
rect 10 -42 14 -32
<< pdcontact >>
rect -10 42 -6 62
rect 0 42 4 62
rect 10 42 14 62
rect -30 5 -26 25
rect -20 5 -16 25
rect -10 5 -6 25
rect 0 5 4 25
rect 10 5 14 25
<< m2contact >>
rect -32 65 -28 69
rect -15 42 -11 62
rect 15 42 19 62
rect -32 28 -28 32
rect 23 -2 27 2
rect -35 -15 -31 -5
rect -43 -22 -39 -18
rect 15 -29 19 -25
rect -15 -42 -11 -32
rect 15 -42 19 -32
rect -35 -49 -31 -45
<< psubstratepcontact >>
rect -26 -44 -22 -36
<< nsubstratencontact >>
rect -25 56 -21 64
<< labels >>
rlabel metal1 -28 65 33 69 1 Vdd
rlabel metal2 -43 -18 -39 75 1 B
rlabel metal1 -31 -49 33 -45 1 Gnd
rlabel metal1 22 35 26 46 1 AddIn
rlabel metal1 -51 42 -15 46 1 AddOut
rlabel metal2 23 -49 27 -2 1 BxnorAdd
<< end >>
