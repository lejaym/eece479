magic
tech scmos
timestamp 1427777783
<< pwell >>
rect 0 395 110 447
rect 0 183 110 284
rect 0 0 110 52
<< nwell >>
rect 0 284 110 395
rect 0 52 110 183
<< polysilicon >>
rect 63 428 84 430
rect 94 428 96 430
rect 16 417 18 419
rect 26 416 48 418
rect 58 416 60 418
rect 16 404 18 407
rect 16 398 22 404
rect 19 384 22 398
rect 26 397 30 416
rect 34 410 48 412
rect 58 410 60 412
rect 16 381 22 384
rect 16 378 18 381
rect 16 356 18 358
rect 26 355 30 391
rect 34 373 37 410
rect 63 393 69 428
rect 72 412 78 419
rect 72 410 84 412
rect 94 410 96 412
rect 72 401 78 410
rect 72 395 94 401
rect 63 373 69 387
rect 89 388 94 395
rect 89 382 105 388
rect 34 371 39 373
rect 59 371 61 373
rect 63 371 74 373
rect 94 371 96 373
rect 63 355 69 371
rect 99 362 105 382
rect 26 353 39 355
rect 59 353 61 355
rect 63 353 74 355
rect 94 353 96 355
rect 26 322 39 324
rect 59 322 61 324
rect 63 322 74 324
rect 94 322 96 324
rect 16 319 18 321
rect 16 296 18 299
rect 16 293 22 296
rect 19 279 22 293
rect 26 286 30 322
rect 63 306 69 322
rect 34 304 39 306
rect 59 304 61 306
rect 63 304 74 306
rect 94 304 96 306
rect 16 273 22 279
rect 16 270 18 273
rect 26 261 30 280
rect 34 267 37 304
rect 63 290 69 304
rect 99 295 105 315
rect 34 265 48 267
rect 58 265 60 267
rect 16 258 18 260
rect 26 259 48 261
rect 58 259 60 261
rect 63 249 69 284
rect 72 289 105 295
rect 72 267 78 289
rect 72 265 84 267
rect 94 265 96 267
rect 72 258 78 265
rect 63 247 84 249
rect 94 247 96 249
rect 39 218 41 220
rect 67 218 69 220
rect 39 206 41 208
rect 67 206 69 208
rect 0 198 28 206
rect 39 202 61 206
rect 67 202 110 206
rect 39 198 41 200
rect 21 186 28 198
rect 56 188 61 202
rect 67 198 69 200
rect 85 198 110 202
rect 39 186 41 188
rect 21 185 53 186
rect 21 179 41 185
rect 21 178 53 179
rect 39 176 41 178
rect 60 176 61 188
rect 67 186 69 188
rect 67 180 77 186
rect 67 176 69 180
rect 39 154 41 156
rect 56 152 61 176
rect 67 154 69 156
rect 85 152 90 198
rect 39 149 61 152
rect 67 149 90 152
rect 39 147 41 149
rect 67 147 69 149
rect 39 125 41 127
rect 67 125 69 127
rect 14 92 28 94
rect 48 92 50 94
rect 53 92 63 94
rect 83 92 85 94
rect 14 31 18 92
rect 53 76 58 92
rect 22 74 28 76
rect 48 74 50 76
rect 53 74 63 76
rect 83 74 85 76
rect 22 37 26 74
rect 53 60 58 74
rect 88 66 94 85
rect 22 35 37 37
rect 47 35 49 37
rect 14 29 37 31
rect 47 29 49 31
rect 53 19 58 54
rect 62 60 94 66
rect 62 37 68 60
rect 62 35 73 37
rect 83 35 85 37
rect 62 28 68 35
rect 53 17 73 19
rect 83 17 85 19
<< ndiffusion >>
rect 84 430 94 431
rect 48 418 58 419
rect 15 407 16 417
rect 18 407 19 417
rect 48 412 58 416
rect 48 409 58 410
rect 84 427 94 428
rect 84 412 94 413
rect 84 409 94 410
rect 15 260 16 270
rect 18 260 19 270
rect 48 267 58 268
rect 48 261 58 265
rect 48 258 58 259
rect 84 267 94 268
rect 84 264 94 265
rect 84 249 94 250
rect 84 246 94 247
rect 38 208 39 218
rect 41 208 42 218
rect 66 208 67 218
rect 69 208 70 218
rect 38 188 39 198
rect 41 188 42 198
rect 66 188 67 198
rect 69 188 70 198
rect 37 37 47 38
rect 37 31 47 35
rect 37 28 47 29
rect 73 37 83 38
rect 73 34 83 35
rect 73 19 83 20
rect 73 16 83 17
<< pdiffusion >>
rect 15 358 16 378
rect 18 358 19 378
rect 39 373 59 374
rect 74 373 94 374
rect 39 370 59 371
rect 39 355 59 356
rect 74 370 94 371
rect 74 355 94 356
rect 39 352 59 353
rect 74 352 94 353
rect 39 324 59 325
rect 74 324 94 325
rect 15 299 16 319
rect 18 299 19 319
rect 39 321 59 322
rect 39 306 59 307
rect 74 321 94 322
rect 74 306 94 307
rect 39 303 59 304
rect 74 303 94 304
rect 38 156 39 176
rect 41 156 42 176
rect 66 156 67 176
rect 69 156 70 176
rect 38 127 39 147
rect 41 127 42 147
rect 66 127 67 147
rect 69 127 70 147
rect 28 94 48 95
rect 63 94 83 95
rect 28 91 48 92
rect 28 76 48 77
rect 63 91 83 92
rect 63 76 83 77
rect 28 73 48 74
rect 63 73 83 74
<< metal1 >>
rect 0 445 110 447
rect 0 441 28 445
rect 35 441 49 445
rect 56 441 71 445
rect 78 441 110 445
rect 0 439 110 441
rect 10 417 15 439
rect 48 423 58 439
rect 84 435 94 439
rect 78 423 84 425
rect 78 420 94 423
rect 10 407 11 417
rect 23 407 31 417
rect 94 413 105 417
rect 10 392 16 398
rect 25 397 31 407
rect 39 391 45 396
rect 25 385 31 391
rect 43 385 45 391
rect 48 393 58 405
rect 74 405 84 409
rect 48 387 63 393
rect 74 391 94 405
rect 98 399 105 413
rect 48 385 69 387
rect 19 381 31 385
rect 19 378 23 381
rect 30 374 39 378
rect 11 346 15 358
rect 30 352 36 374
rect 63 366 69 385
rect 80 383 94 391
rect 74 378 94 383
rect 98 370 105 391
rect 94 366 105 370
rect 39 360 69 366
rect 94 356 99 360
rect 30 348 39 352
rect 30 346 59 348
rect 74 346 94 348
rect 0 344 110 346
rect 0 333 17 344
rect 24 333 42 344
rect 49 333 80 344
rect 87 333 110 344
rect 0 331 110 333
rect 11 319 15 331
rect 30 329 59 331
rect 30 325 39 329
rect 74 329 94 331
rect 30 303 36 325
rect 94 317 99 321
rect 39 311 69 317
rect 30 299 39 303
rect 19 296 23 299
rect 19 292 31 296
rect 63 292 69 311
rect 94 307 105 311
rect 10 279 16 285
rect 25 286 31 292
rect 43 286 45 292
rect 25 270 31 280
rect 39 281 45 286
rect 48 290 69 292
rect 48 284 63 290
rect 74 286 94 299
rect 98 286 105 307
rect 10 260 11 270
rect 23 260 31 270
rect 48 272 58 284
rect 74 278 84 286
rect 92 278 94 286
rect 74 272 94 278
rect 74 268 84 272
rect 98 264 105 278
rect 94 260 105 264
rect 10 238 15 260
rect 48 238 58 254
rect 78 254 94 257
rect 78 252 84 254
rect 84 238 94 242
rect 0 236 110 238
rect 0 224 14 236
rect 21 224 42 236
rect 49 224 71 236
rect 78 224 110 236
rect 0 222 110 224
rect 42 218 46 222
rect 70 218 74 222
rect 10 208 34 218
rect 10 186 20 208
rect 42 198 46 208
rect 0 180 20 186
rect 10 147 20 180
rect 24 185 34 198
rect 49 208 62 218
rect 49 185 53 208
rect 70 198 74 208
rect 58 188 62 198
rect 24 179 29 185
rect 24 156 34 179
rect 42 147 46 156
rect 10 137 34 147
rect 10 131 18 137
rect 24 131 34 137
rect 10 127 34 131
rect 49 147 53 179
rect 60 176 62 188
rect 82 180 110 186
rect 58 156 62 176
rect 70 147 74 156
rect 49 127 62 147
rect 42 123 46 127
rect 70 123 74 127
rect 0 121 110 123
rect 0 110 16 121
rect 23 110 41 121
rect 48 110 79 121
rect 86 110 110 121
rect 0 107 110 110
rect 17 99 23 107
rect 63 99 83 107
rect 17 95 28 99
rect 17 73 23 95
rect 83 87 88 91
rect 28 81 58 87
rect 17 69 28 73
rect 52 64 58 81
rect 83 77 101 81
rect 28 51 34 56
rect 32 45 34 51
rect 37 60 58 64
rect 37 54 52 60
rect 37 42 47 54
rect 50 44 58 54
rect 63 57 83 69
rect 63 49 72 57
rect 80 49 83 57
rect 63 42 83 49
rect 63 38 73 42
rect 88 50 101 77
rect 88 42 92 50
rect 100 42 101 50
rect 88 34 101 42
rect 83 30 101 34
rect 14 17 20 23
rect 37 8 47 24
rect 68 24 83 27
rect 68 22 73 24
rect 73 8 83 12
rect 0 6 110 8
rect 0 2 28 6
rect 35 2 65 6
rect 72 2 86 6
rect 93 2 110 6
rect 0 0 110 2
<< metal2 >>
rect 9 407 60 415
rect 9 392 18 407
rect 9 386 10 392
rect 16 386 18 392
rect 36 396 39 402
rect 45 396 46 402
rect 36 368 46 396
rect 16 359 46 368
rect 16 294 24 359
rect 52 339 60 407
rect 72 391 80 447
rect 10 291 24 294
rect 16 285 24 291
rect 10 283 24 285
rect 16 137 24 283
rect 16 131 18 137
rect 16 20 24 131
rect 29 332 60 339
rect 29 283 37 332
rect 84 286 92 447
rect 29 281 45 283
rect 29 275 39 281
rect 96 391 97 399
rect 96 286 105 391
rect 96 278 97 286
rect 29 273 45 275
rect 29 185 37 273
rect 35 179 37 185
rect 29 62 37 179
rect 34 56 37 62
rect 28 55 37 56
rect 14 17 24 20
rect 20 11 24 17
rect 57 49 72 57
rect 96 50 105 278
rect 57 0 65 49
rect 100 42 105 50
rect 96 0 105 42
<< ntransistor >>
rect 84 428 94 430
rect 16 407 18 417
rect 48 416 58 418
rect 48 410 58 412
rect 84 410 94 412
rect 16 260 18 270
rect 48 265 58 267
rect 48 259 58 261
rect 84 265 94 267
rect 84 247 94 249
rect 39 208 41 218
rect 67 208 69 218
rect 39 188 41 198
rect 67 188 69 198
rect 37 35 47 37
rect 37 29 47 31
rect 73 35 83 37
rect 73 17 83 19
<< ptransistor >>
rect 16 358 18 378
rect 39 371 59 373
rect 74 371 94 373
rect 39 353 59 355
rect 74 353 94 355
rect 39 322 59 324
rect 74 322 94 324
rect 16 299 18 319
rect 39 304 59 306
rect 74 304 94 306
rect 39 156 41 176
rect 67 156 69 176
rect 39 127 41 147
rect 67 127 69 147
rect 28 92 48 94
rect 63 92 83 94
rect 28 74 48 76
rect 63 74 83 76
<< polycontact >>
rect 10 398 16 404
rect 25 391 31 397
rect 72 419 78 425
rect 37 385 43 391
rect 63 387 69 393
rect 99 356 105 362
rect 99 315 105 321
rect 25 280 31 286
rect 10 273 16 279
rect 37 286 43 292
rect 63 284 69 290
rect 72 252 78 258
rect 41 179 53 185
rect 56 176 60 188
rect 77 180 82 186
rect 88 85 94 91
rect 52 54 58 60
rect 26 45 32 51
rect 14 23 20 29
rect 62 22 68 28
<< ndcontact >>
rect 84 431 94 435
rect 48 419 58 423
rect 11 407 15 417
rect 19 407 23 417
rect 48 405 58 409
rect 84 423 94 427
rect 84 413 94 417
rect 84 405 94 409
rect 11 260 15 270
rect 19 260 23 270
rect 48 268 58 272
rect 48 254 58 258
rect 84 268 94 272
rect 84 260 94 264
rect 84 250 94 254
rect 84 242 94 246
rect 34 208 38 218
rect 42 208 46 218
rect 62 208 66 218
rect 70 208 74 218
rect 34 188 38 198
rect 42 188 46 198
rect 62 188 66 198
rect 70 188 74 198
rect 37 38 47 42
rect 37 24 47 28
rect 73 38 83 42
rect 73 30 83 34
rect 73 20 83 24
rect 73 12 83 16
<< pdcontact >>
rect 11 358 15 378
rect 19 358 23 378
rect 39 374 59 378
rect 74 374 94 378
rect 39 366 59 370
rect 39 356 59 360
rect 74 366 94 370
rect 74 356 94 360
rect 39 348 59 352
rect 74 348 94 352
rect 39 325 59 329
rect 74 325 94 329
rect 11 299 15 319
rect 19 299 23 319
rect 39 317 59 321
rect 39 307 59 311
rect 74 317 94 321
rect 74 307 94 311
rect 39 299 59 303
rect 74 299 94 303
rect 34 156 38 176
rect 42 156 46 176
rect 62 156 66 176
rect 70 156 74 176
rect 34 127 38 147
rect 42 127 46 147
rect 62 127 66 147
rect 70 127 74 147
rect 28 95 48 99
rect 63 95 83 99
rect 28 87 48 91
rect 28 77 48 81
rect 63 87 83 91
rect 63 77 83 81
rect 28 69 48 73
rect 63 69 83 73
<< m2contact >>
rect 10 386 16 392
rect 39 396 45 402
rect 97 391 105 399
rect 72 383 80 391
rect 10 285 16 291
rect 39 275 45 281
rect 84 278 92 286
rect 97 278 105 286
rect 29 179 35 185
rect 18 131 24 137
rect 28 56 34 62
rect 72 49 80 57
rect 92 42 100 50
rect 14 11 20 17
<< psubstratepcontact >>
rect 28 441 35 445
rect 49 441 56 445
rect 71 441 78 445
rect 14 224 21 236
rect 42 224 49 236
rect 71 224 78 236
rect 28 2 35 6
rect 65 2 72 6
rect 86 2 93 6
<< nsubstratencontact >>
rect 17 333 24 344
rect 42 333 49 344
rect 80 333 87 344
rect 16 110 23 121
rect 41 110 48 121
rect 79 110 86 121
<< labels >>
rlabel metal1 82 181 97 185 0 S1
rlabel polysilicon 90 198 105 206 0 S0
rlabel metal2 96 115 105 345 0 MUXOUT
rlabel metal2 57 0 65 57 0 REGIN
rlabel metal2 96 50 105 278 0 MUXOUT
rlabel m2contact 84 278 92 286 0 ADDSUB
rlabel m2contact 72 383 80 391 0 DIVIN
rlabel metal1 5 0 28 8 0 GND
rlabel metal1 48 107 79 123 0 Vdd
<< end >>
