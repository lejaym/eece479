magic
tech scmos
timestamp 1427413241
<< pwell >>
rect -30 2 19 38
<< nwell >>
rect -30 -59 19 -2
<< polysilicon >>
rect -29 36 -9 38
rect -29 35 -25 36
rect -11 33 -9 36
rect -1 33 1 35
rect 9 33 11 35
rect -11 22 -9 23
rect -1 22 1 23
rect -11 20 1 22
rect -23 16 -19 18
rect -21 15 -19 16
rect -21 -5 -19 5
rect -21 -27 -19 -25
rect -11 -37 -9 20
rect -1 15 1 17
rect 9 15 11 23
rect 9 11 12 15
rect -1 2 1 5
rect -1 -5 1 -2
rect -1 -28 1 -25
rect -1 -37 1 -35
rect 9 -37 11 11
rect -11 -57 -9 -56
rect -1 -57 1 -56
rect -21 -59 1 -57
rect -21 -63 -19 -59
rect 9 -63 11 -56
<< ndiffusion >>
rect -13 23 -11 33
rect -9 23 -7 33
rect -3 23 -1 33
rect 1 23 3 33
rect 7 23 9 33
rect 11 23 13 33
rect -23 5 -21 15
rect -19 5 -17 15
rect -3 5 -1 15
rect 1 5 3 15
<< pdiffusion >>
rect -23 -25 -21 -5
rect -19 -25 -17 -5
rect -3 -25 -1 -5
rect 1 -25 3 -5
rect -13 -56 -11 -37
rect -9 -56 -7 -37
rect -3 -56 -1 -37
rect 1 -56 3 -37
rect 7 -56 9 -37
rect 11 -56 13 -37
<< metal1 >>
rect -34 38 19 42
rect -25 31 -24 35
rect -7 33 -3 38
rect 13 33 15 38
rect -24 22 -20 23
rect -17 15 -13 23
rect 3 15 7 23
rect 12 15 16 16
rect -27 2 -23 5
rect -8 2 -5 5
rect -44 -2 -40 2
rect -27 -2 -5 2
rect 2 -2 20 2
rect -27 -5 -23 -2
rect -8 -5 -5 -2
rect -27 -40 -23 -25
rect -17 -37 -13 -25
rect -4 -32 -3 -28
rect 4 -37 7 -25
rect -27 -44 -24 -40
rect -26 -59 -22 -58
rect -7 -59 -3 -56
rect 13 -59 17 -56
rect -34 -63 19 -59
<< metal2 >>
rect 4 35 8 42
rect -28 31 -24 35
rect -20 31 8 35
rect -20 23 16 27
rect 12 20 16 23
rect -40 -56 -36 -2
rect -32 -32 -8 -28
rect -32 -48 -28 -32
rect -20 -44 2 -40
rect -32 -52 -8 -48
rect -40 -60 -30 -56
rect -34 -63 -30 -60
rect -12 -63 -8 -52
rect -2 -63 2 -44
<< ntransistor >>
rect -11 23 -9 33
rect -1 23 1 33
rect 9 23 11 33
rect -21 5 -19 15
rect -1 5 1 15
<< ptransistor >>
rect -21 -25 -19 -5
rect -1 -25 1 -5
rect -11 -56 -9 -37
rect -1 -56 1 -37
rect 9 -56 11 -37
<< polycontact >>
rect -29 31 -25 35
rect -24 18 -20 22
rect 12 11 16 15
rect -2 -2 2 2
rect -3 -32 1 -28
<< ndcontact >>
rect -17 23 -13 33
rect -7 23 -3 33
rect 3 23 7 33
rect 13 23 17 33
rect -27 5 -23 15
rect -17 5 -13 15
rect -8 5 -3 15
rect 3 5 7 15
<< pdcontact >>
rect -27 -25 -23 -5
rect -17 -25 -13 -5
rect -8 -25 -3 -5
rect 3 -25 7 -5
rect -17 -56 -13 -37
rect -7 -56 -3 -37
rect 3 -56 7 -37
rect 13 -56 17 -37
<< m2contact >>
rect -24 31 -20 35
rect -24 23 -20 27
rect 12 16 16 20
rect -40 -2 -36 2
rect -8 -32 -4 -28
rect -24 -44 -20 -40
<< psubstratepcontact >>
rect 15 33 19 38
<< nsubstratencontact >>
rect -26 -58 -22 -53
<< labels >>
rlabel polysilicon -1 -5 1 -2 1 Cin
rlabel metal1 -27 -2 -5 2 1 X
rlabel metal1 -34 38 19 42 5 Gnd
rlabel metal1 -34 -63 19 -59 1 Vdd
rlabel space -32 -66 -28 35 3 BxnorAdd
rlabel metal2 -20 23 16 27 1 A
rlabel metal2 4 31 8 42 1 BxnorAdd
rlabel metal1 -44 -2 -40 2 3 Cout
<< end >>
