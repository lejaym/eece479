magic
tech scmos
timestamp 1427936616
<< pwell >>
rect -16 -23 14 -2
<< nwell >>
rect -16 2 14 33
<< polysilicon >>
rect -7 25 -5 27
rect 3 25 5 27
rect -7 -5 -5 5
rect 3 -5 5 5
rect -7 -23 -5 -15
rect 3 -23 5 -15
<< ndiffusion >>
rect -9 -15 -7 -5
rect -5 -15 -3 -5
rect 1 -15 3 -5
rect 5 -15 7 -5
<< pdiffusion >>
rect -9 5 -7 25
rect -5 5 -3 25
rect 1 5 3 25
rect 5 5 7 25
<< metal1 >>
rect -16 29 -6 33
rect 4 29 14 33
rect -13 25 -9 29
rect 7 2 11 5
rect -16 -2 11 2
rect -3 -5 1 -2
rect -13 -19 -9 -15
rect 7 -19 11 -15
rect -16 -23 -4 -19
rect 2 -23 14 -19
<< ntransistor >>
rect -7 -15 -5 -5
rect 3 -15 5 -5
<< ptransistor >>
rect -7 5 -5 25
rect 3 5 5 25
<< ndcontact >>
rect -13 -15 -9 -5
rect -3 -15 1 -5
rect 7 -15 11 -5
<< pdcontact >>
rect -13 5 -9 25
rect -3 5 1 25
rect 7 5 11 25
<< psubstratepcontact >>
rect -4 -23 2 -19
<< nsubstratencontact >>
rect -6 29 4 33
<< labels >>
rlabel nwell -16 2 14 33 1 Vdd
rlabel polysilicon 3 -5 5 5 1 B
rlabel polysilicon -7 -5 -5 5 1 A
rlabel metal1 -16 -2 11 2 1 Out
rlabel metal1 2 -23 14 -19 1 Gnd
<< end >>
