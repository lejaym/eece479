magic
tech scmos
timestamp 1427941063
<< pwell >>
rect -25 -23 14 -2
<< nwell >>
rect -25 2 14 33
<< polysilicon >>
rect -16 25 -14 27
rect -6 25 -4 27
rect 4 25 6 27
rect -16 2 -14 5
rect -16 -5 -14 -2
rect -6 -5 -4 5
rect 4 -5 6 5
rect -16 -17 -14 -15
rect -6 -23 -4 -15
rect 4 -23 6 -15
<< ndiffusion >>
rect -18 -15 -16 -5
rect -14 -15 -12 -5
rect -8 -15 -6 -5
rect -4 -15 -2 -5
rect 2 -15 4 -5
rect 6 -15 8 -5
<< pdiffusion >>
rect -18 5 -16 25
rect -14 5 -12 25
rect -8 5 -6 25
rect -4 5 -2 25
rect 2 5 4 25
rect 6 5 8 25
<< metal1 >>
rect -25 29 -20 33
rect -10 29 14 33
rect -12 25 -8 29
rect 8 25 12 29
rect -24 5 -22 25
rect -24 2 -20 5
rect -2 2 2 5
rect -25 -2 -20 2
rect -13 -2 12 2
rect -24 -5 -20 -2
rect 8 -5 12 -2
rect -24 -15 -22 -5
rect -12 -19 -8 -15
rect -25 -23 -20 -19
rect -10 -23 14 -19
<< ntransistor >>
rect -16 -15 -14 -5
rect -6 -15 -4 -5
rect 4 -15 6 -5
<< ptransistor >>
rect -16 5 -14 25
rect -6 5 -4 25
rect 4 5 6 25
<< polycontact >>
rect -17 -2 -13 2
<< ndcontact >>
rect -22 -15 -18 -5
rect -12 -15 -8 -5
rect -2 -15 2 -5
rect 8 -15 12 -5
<< pdcontact >>
rect -22 5 -18 25
rect -12 5 -8 25
rect -2 5 2 25
rect 8 5 12 25
<< psubstratepcontact >>
rect -20 -23 -10 -19
<< nsubstratencontact >>
rect -20 29 -10 33
<< labels >>
rlabel polysilicon 4 -23 6 -15 1 B
rlabel polysilicon -6 -23 -4 -15 1 A
rlabel metal1 -10 29 14 33 5 Vdd
rlabel metal1 -10 -23 14 -19 1 Gnd
rlabel metal1 -24 -5 -20 5 3 AandB
<< end >>
