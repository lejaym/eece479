magic
tech scmos
timestamp 1427777669
<< polysilicon >>
rect -28 457 -26 459
rect 65 456 67 458
rect 90 456 92 458
rect -28 445 -26 447
rect -28 437 -26 439
rect 65 427 67 436
rect -28 425 -26 427
rect -28 415 -26 417
rect 76 403 81 441
rect 90 434 92 436
rect 90 431 105 434
rect 90 427 92 429
rect 90 403 92 407
rect 76 397 92 403
rect -28 393 -26 395
rect -28 386 -26 388
rect 76 374 81 397
rect 90 395 92 397
rect 90 383 92 385
rect 100 381 105 431
rect 90 377 105 381
rect 90 375 92 377
rect -28 364 -26 366
rect 100 374 105 377
rect 90 363 92 365
rect 35 341 37 343
rect 81 341 83 343
rect -27 339 -25 341
rect 35 329 37 331
rect 81 329 83 331
rect -27 327 -25 329
rect 35 321 37 323
rect 81 321 83 323
rect -27 319 -25 321
rect 35 309 37 311
rect 81 309 83 311
rect -27 307 -25 309
rect 35 299 37 301
rect 81 299 83 301
rect -27 297 -25 299
rect 35 277 37 279
rect 81 277 83 279
rect -27 275 -25 277
rect 35 270 37 272
rect 81 270 83 272
rect -27 268 -25 270
rect 35 248 37 250
rect 81 248 83 250
rect -27 246 -25 248
rect 30 226 32 228
rect 75 226 77 228
rect 30 204 32 206
rect 11 201 32 204
rect 11 154 22 201
rect 30 197 32 199
rect 30 173 32 177
rect 41 173 47 206
rect 75 204 77 206
rect 30 169 47 173
rect 30 165 32 167
rect 18 151 22 154
rect 30 151 32 155
rect 18 147 32 151
rect 30 145 32 147
rect 41 145 47 169
rect 57 201 77 204
rect 57 152 67 201
rect 75 197 77 199
rect 75 173 77 177
rect 86 173 92 206
rect 75 169 92 173
rect 75 165 77 167
rect 63 151 67 152
rect 75 151 77 155
rect 63 147 77 151
rect 63 146 67 147
rect 75 145 77 147
rect 86 145 92 169
rect 30 133 32 135
rect 75 133 77 135
rect 39 111 41 113
rect 67 111 69 113
rect 39 99 41 101
rect 67 99 69 101
rect 0 91 28 99
rect 39 95 61 99
rect 67 95 110 99
rect 39 91 41 93
rect 21 79 28 91
rect 56 81 61 95
rect 67 91 69 93
rect 85 91 110 95
rect 39 79 41 81
rect 21 78 53 79
rect 21 72 41 78
rect 21 71 53 72
rect 39 69 41 71
rect 60 69 61 81
rect 67 79 69 81
rect 67 73 77 79
rect 67 69 69 73
rect 39 47 41 49
rect 56 45 61 69
rect 67 47 69 49
rect 85 45 90 91
rect 39 42 61 45
rect 67 42 90 45
rect 39 40 41 42
rect 67 40 69 42
rect 39 18 41 20
rect 67 18 69 20
<< ndiffusion >>
rect -29 447 -28 457
rect -26 447 -25 457
rect -29 427 -28 437
rect -26 427 -25 437
rect 89 385 90 395
rect 92 385 93 395
rect 89 365 90 375
rect 92 365 93 375
rect -28 329 -27 339
rect -25 329 -24 339
rect 34 331 35 341
rect 37 331 38 341
rect 80 331 81 341
rect 83 331 84 341
rect -28 309 -27 319
rect -25 309 -24 319
rect 34 311 35 321
rect 37 311 38 321
rect 80 311 81 321
rect 83 311 84 321
rect 29 155 30 165
rect 32 155 33 165
rect 74 155 75 165
rect 77 155 78 165
rect 29 135 30 145
rect 32 135 33 145
rect 74 135 75 145
rect 77 135 78 145
rect 38 101 39 111
rect 41 101 42 111
rect 66 101 67 111
rect 69 101 70 111
rect 38 81 39 91
rect 41 81 42 91
rect 66 81 67 91
rect 69 81 70 91
<< pdiffusion >>
rect 64 436 65 456
rect 67 436 68 456
rect -29 395 -28 415
rect -26 395 -25 415
rect 89 436 90 456
rect 92 436 93 456
rect 89 407 90 427
rect 92 407 93 427
rect -29 366 -28 386
rect -26 366 -25 386
rect -28 277 -27 297
rect -25 277 -24 297
rect 34 279 35 299
rect 37 279 38 299
rect 80 279 81 299
rect 83 279 84 299
rect -28 248 -27 268
rect -25 248 -24 268
rect 34 250 35 270
rect 37 250 38 270
rect 80 250 81 270
rect 83 250 84 270
rect 29 206 30 226
rect 32 206 33 226
rect 74 206 75 226
rect 77 206 78 226
rect 29 177 30 197
rect 32 177 33 197
rect 74 177 75 197
rect 77 177 78 197
rect 38 49 39 69
rect 41 49 42 69
rect 66 49 67 69
rect 69 49 70 69
rect 38 20 39 40
rect 41 20 42 40
rect 66 20 67 40
rect 69 20 70 40
<< metal1 >>
rect 0 473 110 476
rect 0 462 16 473
rect 23 462 41 473
rect 48 462 79 473
rect 86 462 110 473
rect 0 460 110 462
rect 68 456 72 460
rect 93 456 97 460
rect 76 452 85 456
rect 81 441 85 452
rect 76 436 85 441
rect 93 427 97 436
rect 70 421 85 427
rect 64 417 85 421
rect 79 385 85 417
rect 64 380 85 385
rect 64 374 69 380
rect 93 375 97 385
rect 0 366 9 374
rect 76 374 85 375
rect 81 366 85 374
rect 76 365 85 366
rect 106 366 110 374
rect 93 361 97 365
rect 0 359 110 361
rect 0 347 14 359
rect 21 347 42 359
rect 49 347 83 359
rect 90 347 110 359
rect 0 345 110 347
rect 0 244 110 246
rect 0 232 16 244
rect 23 232 41 244
rect 48 232 79 244
rect 86 232 110 244
rect 0 230 110 232
rect 25 226 29 230
rect 70 226 74 230
rect 13 197 20 213
rect 37 212 47 226
rect 37 206 41 212
rect 82 212 92 226
rect 82 206 86 212
rect 13 177 25 197
rect 37 177 70 197
rect 82 177 100 197
rect 13 176 29 177
rect 22 165 29 176
rect 37 165 74 177
rect 88 165 100 177
rect 22 155 25 165
rect 37 155 70 165
rect 82 155 100 165
rect 11 143 18 147
rect 11 137 15 143
rect 37 139 41 145
rect 37 135 47 139
rect 57 141 63 146
rect 82 139 86 145
rect 82 135 92 139
rect 25 131 29 135
rect 70 131 74 135
rect 0 129 110 131
rect 0 117 14 129
rect 21 117 42 129
rect 49 117 71 129
rect 78 117 110 129
rect 0 115 110 117
rect 42 111 46 115
rect 70 111 74 115
rect 10 109 34 111
rect 10 103 18 109
rect 24 103 34 109
rect 10 101 34 103
rect 10 79 20 101
rect 42 91 46 101
rect 0 73 20 79
rect 10 40 20 73
rect 24 78 34 91
rect 49 101 62 111
rect 49 78 53 101
rect 70 91 74 101
rect 58 81 62 91
rect 24 72 29 78
rect 24 49 34 72
rect 42 40 46 49
rect 10 20 34 40
rect 49 40 53 72
rect 60 69 62 81
rect 82 73 110 79
rect 58 49 62 69
rect 70 40 74 49
rect 49 20 62 40
rect 42 16 46 20
rect 70 16 74 20
rect 0 14 110 16
rect 0 3 16 14
rect 23 3 41 14
rect 48 3 79 14
rect 86 3 110 14
rect 0 0 110 3
<< metal2 >>
rect 15 143 24 145
rect 21 137 24 143
rect 15 109 24 137
rect 15 103 18 109
rect 15 102 24 103
rect 35 72 37 78
<< ntransistor >>
rect -28 447 -26 457
rect -28 427 -26 437
rect 90 385 92 395
rect 90 365 92 375
rect -27 329 -25 339
rect 35 331 37 341
rect 81 331 83 341
rect -27 309 -25 319
rect 35 311 37 321
rect 81 311 83 321
rect 30 155 32 165
rect 75 155 77 165
rect 30 135 32 145
rect 75 135 77 145
rect 39 101 41 111
rect 67 101 69 111
rect 39 81 41 91
rect 67 81 69 91
<< ptransistor >>
rect 65 436 67 456
rect -28 395 -26 415
rect 90 436 92 456
rect 90 407 92 427
rect -28 366 -26 386
rect -27 277 -25 297
rect 35 279 37 299
rect 81 279 83 299
rect -27 248 -25 268
rect 35 250 37 270
rect 81 250 83 270
rect 30 206 32 226
rect 75 206 77 226
rect 30 177 32 197
rect 75 177 77 197
rect 39 49 41 69
rect 67 49 69 69
rect 39 20 41 40
rect 67 20 69 40
<< polycontact >>
rect 76 441 81 452
rect 64 421 70 427
rect 76 366 81 374
rect 100 366 106 374
rect 41 206 47 212
rect 86 206 92 212
rect 11 147 18 154
rect 57 146 63 152
rect 41 139 47 145
rect 86 139 92 145
rect 41 72 53 78
rect 56 69 60 81
rect 77 73 82 79
<< ndcontact >>
rect -33 447 -29 457
rect -25 447 -21 457
rect -33 427 -29 437
rect -25 427 -21 437
rect 85 385 89 395
rect 93 385 97 395
rect 85 365 89 375
rect 93 365 97 375
rect -32 329 -28 339
rect -24 329 -20 339
rect 30 331 34 341
rect 38 331 42 341
rect 76 331 80 341
rect 84 331 88 341
rect -32 309 -28 319
rect -24 309 -20 319
rect 30 311 34 321
rect 38 311 42 321
rect 76 311 80 321
rect 84 311 88 321
rect 25 155 29 165
rect 33 155 37 165
rect 70 155 74 165
rect 78 155 82 165
rect 25 135 29 145
rect 33 135 37 145
rect 70 135 74 145
rect 78 135 82 145
rect 34 101 38 111
rect 42 101 46 111
rect 62 101 66 111
rect 70 101 74 111
rect 34 81 38 91
rect 42 81 46 91
rect 62 81 66 91
rect 70 81 74 91
<< pdcontact >>
rect 60 436 64 456
rect 68 436 72 456
rect -33 395 -29 415
rect -25 395 -21 415
rect 85 436 89 456
rect 93 436 97 456
rect 85 407 89 427
rect 93 407 97 427
rect -33 366 -29 386
rect -25 366 -21 386
rect -32 277 -28 297
rect -24 277 -20 297
rect 30 279 34 299
rect 38 279 42 299
rect 76 279 80 299
rect 84 279 88 299
rect -32 248 -28 268
rect -24 248 -20 268
rect 30 250 34 270
rect 38 250 42 270
rect 76 250 80 270
rect 84 250 88 270
rect 25 206 29 226
rect 33 206 37 226
rect 70 206 74 226
rect 78 206 82 226
rect 25 177 29 197
rect 33 177 37 197
rect 70 177 74 197
rect 78 177 82 197
rect 34 49 38 69
rect 42 49 46 69
rect 62 49 66 69
rect 70 49 74 69
rect 34 20 38 40
rect 42 20 46 40
rect 62 20 66 40
rect 70 20 74 40
<< m2contact >>
rect 9 366 14 374
rect 64 366 69 374
rect 15 137 21 143
rect 57 135 63 141
rect 18 103 24 109
rect 29 72 35 78
<< psubstratepcontact >>
rect 14 347 21 359
rect 42 347 49 359
rect 83 347 90 359
rect 14 117 21 129
rect 42 117 49 129
rect 71 117 78 129
<< nsubstratencontact >>
rect 16 462 23 473
rect 41 462 48 473
rect 79 462 86 473
rect 16 232 23 244
rect 41 232 48 244
rect 79 232 86 244
rect 16 3 23 14
rect 41 3 48 14
rect 79 3 86 14
<< labels >>
rlabel polysilicon 85 91 105 99 0 CLK
rlabel polysilicon 0 91 28 99 0 INCLK
rlabel metal1 82 73 110 79 0 CLKLD
rlabel metal1 0 73 20 79 0 INCLKCLD
rlabel polysilicon 100 377 105 397 0 RST
<< end >>
