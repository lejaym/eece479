magic
tech scmos
timestamp 1427695733
<< pwell >>
rect 0 68 422 115
<< nwell >>
rect 0 0 422 68
<< polysilicon >>
rect 364 103 366 105
rect 392 103 394 105
rect 32 96 34 98
rect 44 96 65 98
rect 136 96 138 98
rect 148 96 169 98
rect 249 96 251 98
rect 261 96 282 98
rect 23 80 29 89
rect 23 78 34 80
rect 44 78 46 80
rect 13 14 20 34
rect 23 30 29 78
rect 59 61 65 96
rect 68 84 70 86
rect 80 84 103 86
rect 68 78 70 80
rect 80 78 95 80
rect 59 41 65 55
rect 91 41 95 78
rect 32 39 34 41
rect 54 39 65 41
rect 67 39 69 41
rect 89 39 95 41
rect 59 23 65 39
rect 99 23 103 84
rect 127 80 133 89
rect 127 78 138 80
rect 148 78 150 80
rect 127 30 133 78
rect 163 61 169 96
rect 172 84 174 86
rect 184 84 207 86
rect 214 85 216 87
rect 172 78 174 80
rect 184 78 199 80
rect 163 41 169 55
rect 195 41 199 78
rect 136 39 138 41
rect 158 39 169 41
rect 171 39 173 41
rect 193 39 199 41
rect 203 64 207 84
rect 240 80 246 89
rect 240 78 251 80
rect 261 78 263 80
rect 203 58 205 64
rect 163 23 169 39
rect 203 23 207 58
rect 214 46 216 75
rect 240 30 246 78
rect 276 61 282 96
rect 364 91 366 93
rect 392 91 394 93
rect 364 87 386 91
rect 392 87 415 91
rect 285 84 287 86
rect 297 84 320 86
rect 327 85 329 87
rect 285 78 287 80
rect 297 78 312 80
rect 276 41 282 55
rect 308 41 312 78
rect 249 39 251 41
rect 271 39 282 41
rect 284 39 286 41
rect 306 39 312 41
rect 316 64 320 84
rect 364 83 366 85
rect 316 58 318 64
rect 214 24 216 26
rect 276 23 282 39
rect 316 23 320 58
rect 327 46 329 75
rect 381 73 386 87
rect 392 83 394 85
rect 410 81 415 87
rect 364 71 366 73
rect 364 70 378 71
rect 364 66 366 70
rect 364 65 378 66
rect 364 61 366 65
rect 385 61 386 73
rect 392 71 394 73
rect 392 65 402 71
rect 392 61 394 65
rect 364 39 366 41
rect 381 37 386 61
rect 392 39 394 41
rect 410 37 415 75
rect 364 34 386 37
rect 392 34 415 37
rect 364 32 366 34
rect 392 32 394 34
rect 327 24 329 26
rect 32 21 34 23
rect 54 21 65 23
rect 67 21 69 23
rect 89 21 103 23
rect 136 21 138 23
rect 158 21 169 23
rect 171 21 173 23
rect 193 21 207 23
rect 249 21 251 23
rect 271 21 282 23
rect 284 21 286 23
rect 306 21 320 23
rect 13 11 113 14
rect 13 10 122 11
rect 364 10 366 12
rect 392 10 394 12
<< ndiffusion >>
rect 34 98 44 99
rect 138 98 148 99
rect 251 98 261 99
rect 34 95 44 96
rect 34 80 44 81
rect 34 77 44 78
rect 138 95 148 96
rect 70 86 80 87
rect 70 80 80 84
rect 70 77 80 78
rect 138 80 148 81
rect 138 77 148 78
rect 251 95 261 96
rect 174 86 184 87
rect 174 80 184 84
rect 174 77 184 78
rect 213 75 214 85
rect 216 75 217 85
rect 251 80 261 81
rect 251 77 261 78
rect 363 93 364 103
rect 366 93 367 103
rect 391 93 392 103
rect 394 93 395 103
rect 287 86 297 87
rect 287 80 297 84
rect 287 77 297 78
rect 326 75 327 85
rect 329 75 330 85
rect 363 73 364 83
rect 366 73 367 83
rect 391 73 392 83
rect 394 73 395 83
<< pdiffusion >>
rect 34 41 54 42
rect 69 41 89 42
rect 34 38 54 39
rect 34 23 54 24
rect 69 38 89 39
rect 69 23 89 24
rect 138 41 158 42
rect 173 41 193 42
rect 138 38 158 39
rect 138 23 158 24
rect 173 38 193 39
rect 173 23 193 24
rect 213 26 214 46
rect 216 26 217 46
rect 251 41 271 42
rect 286 41 306 42
rect 251 38 271 39
rect 251 23 271 24
rect 286 38 306 39
rect 286 23 306 24
rect 326 26 327 46
rect 329 26 330 46
rect 363 41 364 61
rect 366 41 367 61
rect 391 41 392 61
rect 394 41 395 61
rect 34 20 54 21
rect 69 20 89 21
rect 138 20 158 21
rect 173 20 193 21
rect 251 20 271 21
rect 286 20 306 21
rect 363 12 364 32
rect 366 12 367 32
rect 391 12 392 32
rect 394 12 395 32
<< metal1 >>
rect 0 113 422 115
rect 0 109 45 113
rect 52 109 82 113
rect 89 109 126 113
rect 133 109 165 113
rect 172 109 209 113
rect 216 109 267 113
rect 274 109 315 113
rect 322 109 353 113
rect 360 109 385 113
rect 392 109 422 113
rect 0 107 422 109
rect 34 103 44 107
rect 29 91 34 95
rect 70 91 80 107
rect 138 103 148 107
rect 133 91 138 95
rect 174 91 184 107
rect 217 85 222 107
rect 251 103 261 107
rect 246 91 251 95
rect 287 91 297 107
rect 330 85 335 107
rect 367 103 371 107
rect 395 103 399 107
rect 0 74 7 80
rect 13 81 34 85
rect 117 81 138 85
rect 0 62 7 65
rect 13 41 26 81
rect 44 73 54 77
rect 34 67 54 73
rect 45 49 54 67
rect 34 46 54 49
rect 59 61 67 71
rect 70 61 80 73
rect 65 55 80 61
rect 59 53 80 55
rect 83 64 85 70
rect 83 59 89 64
rect 105 59 111 65
rect 109 53 111 59
rect 59 51 67 53
rect 20 38 26 41
rect 20 34 34 38
rect 59 34 65 51
rect 89 42 100 46
rect 117 42 130 81
rect 153 73 161 77
rect 138 70 161 73
rect 138 67 158 70
rect 149 52 158 67
rect 174 61 184 73
rect 221 75 222 85
rect 230 81 251 85
rect 138 46 158 52
rect 169 55 184 61
rect 163 53 184 55
rect 187 64 189 70
rect 209 68 213 75
rect 204 64 213 68
rect 187 59 193 64
rect 204 58 205 64
rect 211 58 213 64
rect 218 59 224 65
rect 204 54 213 58
rect 59 28 89 34
rect 29 24 34 28
rect 94 20 100 42
rect 89 16 100 20
rect 34 8 54 16
rect 94 8 100 16
rect 113 34 117 42
rect 125 38 130 42
rect 125 34 138 38
rect 163 34 169 53
rect 209 46 213 54
rect 222 53 224 59
rect 193 42 204 46
rect 113 17 122 34
rect 163 28 193 34
rect 133 24 138 28
rect 198 20 204 42
rect 230 42 243 81
rect 266 73 274 77
rect 251 67 271 73
rect 262 52 271 67
rect 287 61 297 73
rect 334 75 335 85
rect 342 93 359 103
rect 251 46 271 52
rect 282 55 297 61
rect 276 53 297 55
rect 322 68 326 75
rect 300 59 306 64
rect 317 64 326 68
rect 335 65 337 71
rect 300 53 302 59
rect 317 58 318 64
rect 324 58 326 64
rect 317 54 326 58
rect 238 38 243 42
rect 238 34 251 38
rect 276 34 282 53
rect 322 46 326 54
rect 331 59 337 65
rect 342 59 348 93
rect 367 83 371 93
rect 306 42 317 46
rect 193 16 204 20
rect 138 8 158 16
rect 198 8 204 16
rect 217 8 221 26
rect 276 28 306 34
rect 246 24 251 28
rect 311 20 317 42
rect 306 16 317 20
rect 251 8 271 16
rect 311 8 317 16
rect 330 8 334 26
rect 342 32 348 53
rect 353 71 359 83
rect 374 93 387 103
rect 374 70 378 93
rect 395 83 399 93
rect 383 73 387 83
rect 415 75 422 81
rect 353 41 359 65
rect 367 32 371 41
rect 342 12 359 32
rect 374 32 378 66
rect 385 61 387 73
rect 407 65 422 71
rect 383 41 387 61
rect 395 32 399 41
rect 374 12 387 32
rect 367 8 371 12
rect 395 8 399 12
rect 0 6 422 8
rect 0 2 41 6
rect 48 2 74 6
rect 81 2 145 6
rect 152 2 182 6
rect 189 2 212 6
rect 219 2 258 6
rect 265 2 296 6
rect 303 2 321 6
rect 328 2 360 6
rect 367 2 388 6
rect 395 2 422 6
rect 0 0 422 2
<< metal2 >>
rect 0 103 113 110
rect 0 87 7 103
rect 103 73 113 103
rect 153 84 161 96
rect 266 84 274 96
rect 103 71 360 73
rect 7 65 67 71
rect 103 65 105 71
rect 111 65 218 71
rect 224 70 353 71
rect 224 65 300 70
rect 0 62 67 65
rect 306 65 353 70
rect 359 65 360 71
rect 59 59 67 62
rect 19 49 34 55
rect 59 53 83 59
rect 89 53 187 59
rect 193 53 331 59
rect 337 53 342 59
rect 348 53 350 59
rect 59 51 350 53
rect 19 0 29 49
rect 114 42 125 45
rect 114 34 117 42
rect 114 19 125 34
rect 228 42 238 44
rect 228 34 230 42
rect 228 19 238 34
rect 114 9 238 19
rect 167 0 175 9
<< ntransistor >>
rect 34 96 44 98
rect 138 96 148 98
rect 251 96 261 98
rect 34 78 44 80
rect 70 84 80 86
rect 70 78 80 80
rect 138 78 148 80
rect 174 84 184 86
rect 174 78 184 80
rect 214 75 216 85
rect 251 78 261 80
rect 364 93 366 103
rect 392 93 394 103
rect 287 84 297 86
rect 287 78 297 80
rect 327 75 329 85
rect 364 73 366 83
rect 392 73 394 83
<< ptransistor >>
rect 34 39 54 41
rect 69 39 89 41
rect 138 39 158 41
rect 173 39 193 41
rect 214 26 216 46
rect 251 39 271 41
rect 286 39 306 41
rect 327 26 329 46
rect 364 41 366 61
rect 392 41 394 61
rect 34 21 54 23
rect 69 21 89 23
rect 138 21 158 23
rect 173 21 193 23
rect 251 21 271 23
rect 286 21 306 23
rect 364 12 366 32
rect 392 12 394 32
<< polycontact >>
rect 23 89 29 95
rect 13 34 20 41
rect 127 89 133 95
rect 85 64 91 70
rect 59 55 65 61
rect 23 24 29 30
rect 103 53 109 59
rect 240 89 246 95
rect 189 64 195 70
rect 163 55 169 61
rect 205 58 211 64
rect 127 24 133 30
rect 216 53 222 59
rect 276 55 282 61
rect 302 53 308 59
rect 318 58 324 64
rect 240 24 246 30
rect 410 75 415 81
rect 329 65 335 71
rect 366 66 378 70
rect 381 61 385 73
rect 402 65 407 71
rect 113 11 122 17
<< ndcontact >>
rect 34 99 44 103
rect 138 99 148 103
rect 251 99 261 103
rect 34 91 44 95
rect 34 81 44 85
rect 34 73 44 77
rect 70 87 80 91
rect 138 91 148 95
rect 70 73 80 77
rect 138 81 148 85
rect 138 73 148 77
rect 174 87 184 91
rect 251 91 261 95
rect 174 73 184 77
rect 209 75 213 85
rect 217 75 221 85
rect 251 81 261 85
rect 251 73 261 77
rect 359 93 363 103
rect 367 93 371 103
rect 387 93 391 103
rect 395 93 399 103
rect 287 87 297 91
rect 287 73 297 77
rect 322 75 326 85
rect 330 75 334 85
rect 359 73 363 83
rect 367 73 371 83
rect 387 73 391 83
rect 395 73 399 83
<< pdcontact >>
rect 34 42 54 46
rect 69 42 89 46
rect 34 34 54 38
rect 34 24 54 28
rect 69 34 89 38
rect 69 24 89 28
rect 138 42 158 46
rect 173 42 193 46
rect 138 34 158 38
rect 138 24 158 28
rect 173 34 193 38
rect 173 24 193 28
rect 209 26 213 46
rect 217 26 221 46
rect 251 42 271 46
rect 286 42 306 46
rect 251 34 271 38
rect 251 24 271 28
rect 286 34 306 38
rect 286 24 306 28
rect 322 26 326 46
rect 330 26 334 46
rect 359 41 363 61
rect 367 41 371 61
rect 387 41 391 61
rect 395 41 399 61
rect 34 16 54 20
rect 69 16 89 20
rect 138 16 158 20
rect 173 16 193 20
rect 251 16 271 20
rect 286 16 306 20
rect 359 12 363 32
rect 367 12 371 32
rect 387 12 391 32
rect 395 12 399 32
<< m2contact >>
rect 0 80 7 87
rect 0 65 7 71
rect 34 49 45 55
rect 105 65 111 71
rect 83 53 89 59
rect 153 77 161 84
rect 187 53 193 59
rect 218 65 224 71
rect 117 34 125 42
rect 266 77 274 84
rect 300 64 306 70
rect 230 34 238 42
rect 331 53 337 59
rect 342 53 348 59
rect 353 65 359 71
<< psubstratepcontact >>
rect 45 109 52 113
rect 82 109 89 113
rect 126 109 133 113
rect 165 109 172 113
rect 209 109 216 113
rect 267 109 274 113
rect 315 109 322 113
rect 353 109 360 113
rect 385 109 392 113
<< nsubstratencontact >>
rect 41 2 48 6
rect 74 2 81 6
rect 145 2 152 6
rect 182 2 189 6
rect 212 2 219 6
rect 258 2 265 6
rect 296 2 303 6
rect 321 2 328 6
rect 360 2 367 6
rect 388 2 395 6
<< labels >>
rlabel metal1 415 76 422 80 0 S0
rlabel metal1 407 66 422 70 0 S1
rlabel metal2 266 84 274 96 0 ADDSUB
rlabel metal2 114 9 238 19 0 MUXOUT
rlabel metal2 19 0 29 55 0 REGIN
rlabel metal2 153 84 161 96 0 DIVIN
rlabel metal1 0 107 422 115 0 GND
rlabel nwell 0 0 422 8 0 Vdd
<< end >>
