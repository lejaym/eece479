magic
tech scmos
timestamp 1427427203
<< pwell >>
rect -54 -70 24 -29
<< nwell >>
rect -54 -25 24 36
<< polysilicon >>
rect -26 5 -24 52
rect -15 36 -14 39
rect -16 33 -14 36
rect -6 36 -5 39
rect -6 33 -4 36
rect -27 1 -24 5
rect -46 -2 -44 0
rect -36 -2 -34 0
rect -26 -2 -24 1
rect -16 -2 -14 13
rect -6 -2 -4 13
rect 4 -2 6 52
rect 14 33 16 35
rect 14 -17 16 13
rect 14 -21 17 -17
rect -46 -25 -44 -22
rect -46 -32 -44 -29
rect -36 -32 -34 -22
rect -26 -32 -24 -22
rect -16 -32 -14 -22
rect -6 -32 -4 -22
rect 4 -25 6 -22
rect 4 -32 6 -29
rect -46 -44 -44 -42
rect -36 -45 -34 -42
rect -26 -44 -24 -42
rect -36 -49 -35 -45
rect -16 -57 -14 -42
rect -6 -57 -4 -42
rect 4 -44 6 -42
rect 14 -57 16 -21
rect -16 -69 -14 -67
rect -6 -69 -4 -67
rect 14 -69 16 -67
<< ndiffusion >>
rect -48 -42 -46 -32
rect -44 -42 -42 -32
rect -38 -42 -36 -32
rect -34 -42 -32 -32
rect -28 -42 -26 -32
rect -24 -42 -22 -32
rect -18 -42 -16 -32
rect -14 -42 -12 -32
rect -8 -42 -6 -32
rect -4 -42 -2 -32
rect 2 -42 4 -32
rect 6 -42 8 -32
rect -18 -67 -16 -57
rect -14 -67 -12 -57
rect -8 -67 -6 -57
rect -4 -67 -2 -57
rect 12 -67 14 -57
rect 16 -67 18 -57
<< pdiffusion >>
rect -18 13 -16 33
rect -14 13 -12 33
rect -8 13 -6 33
rect -4 13 -2 33
rect 12 13 14 33
rect 16 13 18 33
rect -48 -22 -46 -2
rect -44 -22 -42 -2
rect -38 -22 -36 -2
rect -34 -22 -32 -2
rect -28 -22 -26 -2
rect -24 -22 -22 -2
rect -18 -22 -16 -2
rect -14 -22 -12 -2
rect -8 -22 -6 -2
rect -4 -22 -2 -2
rect 2 -22 4 -2
rect 6 -22 8 -2
<< metal1 >>
rect -57 48 24 52
rect -42 25 -38 48
rect -19 40 -15 41
rect -12 33 -8 48
rect -5 40 -1 41
rect 18 33 22 48
rect -42 -2 -38 12
rect -31 5 -27 16
rect -22 5 -18 13
rect -2 12 2 13
rect 8 5 12 13
rect -22 1 12 5
rect -2 -2 2 1
rect 18 -2 22 13
rect -54 -22 -52 -2
rect 12 -6 22 -2
rect 17 -17 21 -13
rect -54 -32 -50 -22
rect -12 -25 -8 -22
rect -43 -29 -8 -25
rect 8 -29 9 -25
rect -12 -32 -8 -29
rect -54 -42 -52 -32
rect 12 -42 22 -38
rect -54 -43 -50 -42
rect -42 -53 -38 -42
rect -2 -45 2 -42
rect -31 -49 -29 -45
rect -22 -49 12 -45
rect -42 -70 -38 -66
rect -22 -57 -18 -49
rect -2 -57 2 -56
rect 8 -57 12 -49
rect 18 -57 22 -42
rect -12 -70 -8 -67
rect 18 -70 22 -67
rect -55 -74 24 -70
<< metal2 >>
rect -39 12 -35 52
rect -17 45 -13 52
rect -15 41 -13 45
rect -7 45 -3 52
rect -7 41 -5 45
rect -27 16 21 20
rect -39 8 -2 12
rect -54 -74 -50 -47
rect -29 -60 -25 -49
rect -2 -52 2 8
rect 17 -9 21 16
rect 9 -60 13 -29
rect -29 -64 13 -60
<< ntransistor >>
rect -46 -42 -44 -32
rect -36 -42 -34 -32
rect -26 -42 -24 -32
rect -16 -42 -14 -32
rect -6 -42 -4 -32
rect 4 -42 6 -32
rect -16 -67 -14 -57
rect -6 -67 -4 -57
rect 14 -67 16 -57
<< ptransistor >>
rect -16 13 -14 33
rect -6 13 -4 33
rect 14 13 16 33
rect -46 -22 -44 -2
rect -36 -22 -34 -2
rect -26 -22 -24 -2
rect -16 -22 -14 -2
rect -6 -22 -4 -2
rect 4 -22 6 -2
<< polycontact >>
rect -19 36 -15 40
rect -5 36 -1 40
rect -31 1 -27 5
rect 17 -21 21 -17
rect -47 -29 -43 -25
rect 4 -29 8 -25
rect -35 -49 -31 -45
<< ndcontact >>
rect -52 -42 -48 -32
rect -42 -42 -38 -32
rect -32 -42 -28 -32
rect -22 -42 -18 -32
rect -12 -42 -8 -32
rect -2 -42 2 -32
rect 8 -42 12 -32
rect -22 -67 -18 -57
rect -12 -67 -8 -57
rect -2 -67 2 -57
rect 8 -67 12 -57
rect 18 -67 22 -57
<< pdcontact >>
rect -22 13 -18 33
rect -12 13 -8 33
rect -2 13 2 33
rect 8 13 12 33
rect 18 13 22 33
rect -52 -22 -48 -2
rect -42 -22 -38 -2
rect -32 -22 -28 -2
rect -22 -22 -18 -2
rect -12 -22 -8 -2
rect -2 -22 2 -2
rect 8 -22 12 -2
<< m2contact >>
rect -19 41 -15 45
rect -5 41 -1 45
rect -31 16 -27 20
rect -2 8 2 12
rect 17 -13 21 -9
rect 9 -29 13 -25
rect -54 -47 -50 -43
rect -29 -49 -25 -45
rect -2 -56 2 -52
<< psubstratepcontact >>
rect -42 -66 -38 -53
<< nsubstratencontact >>
rect -42 12 -38 25
<< labels >>
rlabel polysilicon 4 -2 6 35 1 A
rlabel metal1 -55 -74 24 -70 1 Gnd
rlabel metal2 -54 -74 -50 -47 3 sum
rlabel metal1 -57 48 24 52 5 Vdd
rlabel metal2 -7 45 -3 52 5 X
rlabel metal2 -17 45 -13 52 5 Cin
rlabel metal2 -39 8 -35 52 1 Cout
rlabel polysilicon -26 -2 -24 52 1 BxnorAdd
<< end >>
