magic
tech scmos
timestamp 1427755732
<< pwell >>
rect 0 280 100 332
rect 0 68 100 169
rect 0 -115 100 -63
<< nwell >>
rect 0 169 100 280
rect 0 -63 100 68
<< polysilicon >>
rect 58 313 79 315
rect 89 313 91 315
rect 11 302 13 304
rect 21 301 43 303
rect 53 301 55 303
rect 11 289 13 292
rect 11 283 17 289
rect 14 270 17 283
rect 21 282 25 301
rect 29 295 43 297
rect 53 295 55 297
rect 21 270 25 276
rect 14 269 25 270
rect 11 266 25 269
rect 11 263 13 266
rect 11 241 13 243
rect 21 240 25 266
rect 29 258 32 295
rect 58 278 64 313
rect 67 297 73 304
rect 67 295 79 297
rect 89 295 91 297
rect 67 286 73 295
rect 67 280 89 286
rect 58 258 64 272
rect 84 273 89 280
rect 84 267 100 273
rect 29 256 34 258
rect 54 256 56 258
rect 58 256 69 258
rect 89 256 91 258
rect 58 240 64 256
rect 94 247 100 267
rect 21 238 34 240
rect 54 238 56 240
rect 58 238 69 240
rect 89 238 91 240
rect 21 207 34 209
rect 54 207 56 209
rect 58 207 69 209
rect 89 207 91 209
rect 11 204 13 206
rect 11 181 13 184
rect 21 181 25 207
rect 58 191 64 207
rect 11 178 25 181
rect 14 177 25 178
rect 14 164 17 177
rect 21 171 25 177
rect 29 189 34 191
rect 54 189 56 191
rect 58 189 69 191
rect 89 189 91 191
rect 11 158 17 164
rect 11 155 13 158
rect 21 146 25 165
rect 29 152 32 189
rect 58 175 64 189
rect 94 180 100 200
rect 29 150 43 152
rect 53 150 55 152
rect 11 143 13 145
rect 21 144 43 146
rect 53 144 55 146
rect 58 134 64 169
rect 67 174 100 180
rect 67 152 73 174
rect 67 150 79 152
rect 89 150 91 152
rect 67 143 73 150
rect 58 132 79 134
rect 89 132 91 134
rect 34 103 36 105
rect 62 103 64 105
rect 34 91 36 93
rect 62 91 64 93
rect 0 83 23 91
rect 34 87 56 91
rect 62 87 100 91
rect 34 83 36 85
rect 16 71 23 83
rect 51 73 56 87
rect 62 83 64 85
rect 80 83 100 87
rect 34 71 36 73
rect 16 70 48 71
rect 16 64 36 70
rect 16 63 48 64
rect 34 61 36 63
rect 55 61 56 73
rect 62 71 64 73
rect 62 65 72 71
rect 62 61 64 65
rect 34 39 36 41
rect 51 37 56 61
rect 62 39 64 41
rect 80 37 85 83
rect 34 34 56 37
rect 62 34 85 37
rect 34 32 36 34
rect 62 32 64 34
rect 34 10 36 12
rect 62 10 64 12
rect 9 -23 23 -21
rect 43 -23 45 -21
rect 48 -23 58 -21
rect 78 -23 80 -21
rect 9 -84 13 -23
rect 48 -39 53 -23
rect 17 -41 23 -39
rect 43 -41 45 -39
rect 48 -41 58 -39
rect 78 -41 80 -39
rect 17 -78 21 -41
rect 48 -55 53 -41
rect 83 -49 89 -30
rect 17 -80 32 -78
rect 42 -80 44 -78
rect 9 -86 32 -84
rect 42 -86 44 -84
rect 48 -96 53 -61
rect 57 -55 89 -49
rect 57 -78 63 -55
rect 57 -80 68 -78
rect 78 -80 80 -78
rect 57 -87 63 -80
rect 48 -98 68 -96
rect 78 -98 80 -96
<< ndiffusion >>
rect 79 315 89 316
rect 43 303 53 304
rect 10 292 11 302
rect 13 292 14 302
rect 43 297 53 301
rect 43 294 53 295
rect 79 312 89 313
rect 79 297 89 298
rect 79 294 89 295
rect 10 145 11 155
rect 13 145 14 155
rect 43 152 53 153
rect 43 146 53 150
rect 43 143 53 144
rect 79 152 89 153
rect 79 149 89 150
rect 79 134 89 135
rect 79 131 89 132
rect 33 93 34 103
rect 36 93 37 103
rect 61 93 62 103
rect 64 93 65 103
rect 33 73 34 83
rect 36 73 37 83
rect 61 73 62 83
rect 64 73 65 83
rect 32 -78 42 -77
rect 32 -84 42 -80
rect 32 -87 42 -86
rect 68 -78 78 -77
rect 68 -81 78 -80
rect 68 -96 78 -95
rect 68 -99 78 -98
<< pdiffusion >>
rect 10 243 11 263
rect 13 243 14 263
rect 34 258 54 259
rect 69 258 89 259
rect 34 255 54 256
rect 34 240 54 241
rect 69 255 89 256
rect 69 240 89 241
rect 34 237 54 238
rect 69 237 89 238
rect 34 209 54 210
rect 69 209 89 210
rect 10 184 11 204
rect 13 184 14 204
rect 34 206 54 207
rect 34 191 54 192
rect 69 206 89 207
rect 69 191 89 192
rect 34 188 54 189
rect 69 188 89 189
rect 33 41 34 61
rect 36 41 37 61
rect 61 41 62 61
rect 64 41 65 61
rect 33 12 34 32
rect 36 12 37 32
rect 61 12 62 32
rect 64 12 65 32
rect 23 -21 43 -20
rect 58 -21 78 -20
rect 23 -24 43 -23
rect 23 -39 43 -38
rect 58 -24 78 -23
rect 58 -39 78 -38
rect 23 -42 43 -41
rect 58 -42 78 -41
<< metal1 >>
rect 110 333 127 334
rect 100 332 127 333
rect 0 330 127 332
rect 0 326 23 330
rect 30 326 44 330
rect 51 326 66 330
rect 73 326 127 330
rect 0 324 127 326
rect 5 302 10 324
rect 43 308 53 324
rect 79 320 89 324
rect 73 308 79 310
rect 73 305 89 308
rect 5 292 6 302
rect 18 292 26 302
rect 89 298 100 302
rect 5 277 11 283
rect 20 282 26 292
rect 34 276 40 281
rect 20 270 26 276
rect 38 270 40 276
rect 43 278 53 290
rect 69 290 79 294
rect 43 272 58 278
rect 69 276 89 290
rect 93 284 100 298
rect 43 270 64 272
rect 14 266 26 270
rect 14 263 18 266
rect 25 259 34 263
rect -26 231 0 232
rect 6 231 10 243
rect 25 237 31 259
rect 58 251 64 270
rect 75 268 89 276
rect 69 263 89 268
rect 93 255 100 276
rect 89 251 100 255
rect 34 245 64 251
rect 89 241 94 245
rect 25 233 34 237
rect 25 231 54 233
rect 69 231 89 233
rect -26 229 100 231
rect -26 218 12 229
rect 19 218 37 229
rect 44 218 75 229
rect 82 218 100 229
rect -27 216 100 218
rect -27 8 -10 216
rect 6 204 10 216
rect 25 214 54 216
rect 25 210 34 214
rect 69 214 89 216
rect 25 188 31 210
rect 89 202 94 206
rect 34 196 64 202
rect 25 184 34 188
rect 14 181 18 184
rect 14 177 26 181
rect 58 177 64 196
rect 89 192 100 196
rect 5 164 11 170
rect 20 171 26 177
rect 38 171 40 177
rect 20 155 26 165
rect 34 166 40 171
rect 43 175 64 177
rect 43 169 58 175
rect 69 171 89 184
rect 93 171 100 192
rect 5 145 6 155
rect 18 145 26 155
rect 43 157 53 169
rect 69 163 79 171
rect 87 163 89 171
rect 69 157 89 163
rect 69 153 79 157
rect 93 149 100 163
rect 89 145 100 149
rect 5 123 10 145
rect 43 123 53 139
rect 73 139 89 142
rect 73 137 79 139
rect 79 123 89 127
rect 110 123 127 324
rect 0 121 127 123
rect 0 109 9 121
rect 16 109 37 121
rect 44 109 66 121
rect 73 111 127 121
rect 73 109 129 111
rect 0 107 129 109
rect 37 103 41 107
rect 65 103 69 107
rect 5 93 29 103
rect 5 71 15 93
rect 37 83 41 93
rect 0 65 15 71
rect 5 32 15 65
rect 19 70 29 83
rect 44 93 57 103
rect 44 70 48 93
rect 65 83 69 93
rect 53 73 57 83
rect 19 64 24 70
rect 19 41 29 64
rect 37 32 41 41
rect 5 22 29 32
rect 5 16 13 22
rect 19 16 29 22
rect 5 12 29 16
rect 44 32 48 64
rect 55 61 57 73
rect 77 65 100 71
rect 53 41 57 61
rect 65 32 69 41
rect 44 12 57 32
rect 37 8 41 12
rect 65 8 69 12
rect -27 6 100 8
rect -27 -5 11 6
rect 18 -5 36 6
rect 43 -5 74 6
rect 81 -5 100 6
rect -27 -8 100 -5
rect 12 -16 18 -8
rect 58 -16 78 -8
rect 12 -20 23 -16
rect 12 -42 18 -20
rect 78 -28 83 -24
rect 23 -34 53 -28
rect 12 -46 23 -42
rect 47 -51 53 -34
rect 78 -38 96 -34
rect 23 -64 29 -59
rect 27 -70 29 -64
rect 32 -55 53 -51
rect 32 -61 47 -55
rect 32 -73 42 -61
rect 45 -71 53 -61
rect 58 -58 78 -46
rect 58 -66 67 -58
rect 75 -66 78 -58
rect 58 -73 78 -66
rect 58 -77 68 -73
rect 83 -65 96 -38
rect 83 -73 87 -65
rect 95 -73 96 -65
rect 83 -81 96 -73
rect 78 -85 96 -81
rect 9 -98 15 -92
rect 32 -107 42 -91
rect 63 -91 78 -88
rect 63 -93 68 -91
rect 68 -107 78 -103
rect 110 -106 129 107
rect 100 -107 129 -106
rect 0 -109 129 -107
rect 0 -113 23 -109
rect 30 -113 60 -109
rect 67 -113 81 -109
rect 88 -113 129 -109
rect 0 -115 129 -113
<< metal2 >>
rect 4 292 55 300
rect 4 277 13 292
rect 4 271 5 277
rect 11 271 13 277
rect 31 281 34 287
rect 40 281 41 287
rect 31 253 41 281
rect 11 244 41 253
rect 11 179 19 244
rect 47 224 55 292
rect 67 276 75 332
rect 5 176 19 179
rect 11 170 19 176
rect 5 168 19 170
rect 11 22 19 168
rect 11 16 13 22
rect 11 -95 19 16
rect 24 217 55 224
rect 24 168 32 217
rect 79 171 87 332
rect 24 166 40 168
rect 24 160 34 166
rect 91 276 92 284
rect 91 171 100 276
rect 91 163 92 171
rect 24 158 40 160
rect 24 70 32 158
rect 30 64 32 70
rect 24 -53 32 64
rect 29 -59 32 -53
rect 23 -60 32 -59
rect 9 -98 19 -95
rect 15 -104 19 -98
rect 52 -66 67 -58
rect 91 -65 100 163
rect 52 -115 60 -66
rect 95 -73 100 -65
rect 91 -115 100 -73
<< ntransistor >>
rect 79 313 89 315
rect 11 292 13 302
rect 43 301 53 303
rect 43 295 53 297
rect 79 295 89 297
rect 11 145 13 155
rect 43 150 53 152
rect 43 144 53 146
rect 79 150 89 152
rect 79 132 89 134
rect 34 93 36 103
rect 62 93 64 103
rect 34 73 36 83
rect 62 73 64 83
rect 32 -80 42 -78
rect 32 -86 42 -84
rect 68 -80 78 -78
rect 68 -98 78 -96
<< ptransistor >>
rect 11 243 13 263
rect 34 256 54 258
rect 69 256 89 258
rect 34 238 54 240
rect 69 238 89 240
rect 34 207 54 209
rect 69 207 89 209
rect 11 184 13 204
rect 34 189 54 191
rect 69 189 89 191
rect 34 41 36 61
rect 62 41 64 61
rect 34 12 36 32
rect 62 12 64 32
rect 23 -23 43 -21
rect 58 -23 78 -21
rect 23 -41 43 -39
rect 58 -41 78 -39
<< polycontact >>
rect 5 283 11 289
rect 20 276 26 282
rect 67 304 73 310
rect 32 270 38 276
rect 58 272 64 278
rect 94 241 100 247
rect 94 200 100 206
rect 20 165 26 171
rect 5 158 11 164
rect 32 171 38 177
rect 58 169 64 175
rect 67 137 73 143
rect 36 64 48 70
rect 51 61 55 73
rect 72 65 77 71
rect 83 -30 89 -24
rect 47 -61 53 -55
rect 21 -70 27 -64
rect 9 -92 15 -86
rect 57 -93 63 -87
<< ndcontact >>
rect 79 316 89 320
rect 43 304 53 308
rect 6 292 10 302
rect 14 292 18 302
rect 43 290 53 294
rect 79 308 89 312
rect 79 298 89 302
rect 79 290 89 294
rect 6 145 10 155
rect 14 145 18 155
rect 43 153 53 157
rect 43 139 53 143
rect 79 153 89 157
rect 79 145 89 149
rect 79 135 89 139
rect 79 127 89 131
rect 29 93 33 103
rect 37 93 41 103
rect 57 93 61 103
rect 65 93 69 103
rect 29 73 33 83
rect 37 73 41 83
rect 57 73 61 83
rect 65 73 69 83
rect 32 -77 42 -73
rect 32 -91 42 -87
rect 68 -77 78 -73
rect 68 -85 78 -81
rect 68 -95 78 -91
rect 68 -103 78 -99
<< pdcontact >>
rect 6 243 10 263
rect 14 243 18 263
rect 34 259 54 263
rect 69 259 89 263
rect 34 251 54 255
rect 34 241 54 245
rect 69 251 89 255
rect 69 241 89 245
rect 34 233 54 237
rect 69 233 89 237
rect 34 210 54 214
rect 69 210 89 214
rect 6 184 10 204
rect 14 184 18 204
rect 34 202 54 206
rect 34 192 54 196
rect 69 202 89 206
rect 69 192 89 196
rect 34 184 54 188
rect 69 184 89 188
rect 29 41 33 61
rect 37 41 41 61
rect 57 41 61 61
rect 65 41 69 61
rect 29 12 33 32
rect 37 12 41 32
rect 57 12 61 32
rect 65 12 69 32
rect 23 -20 43 -16
rect 58 -20 78 -16
rect 23 -28 43 -24
rect 23 -38 43 -34
rect 58 -28 78 -24
rect 58 -38 78 -34
rect 23 -46 43 -42
rect 58 -46 78 -42
<< m2contact >>
rect 5 271 11 277
rect 34 281 40 287
rect 92 276 100 284
rect 67 268 75 276
rect 5 170 11 176
rect 34 160 40 166
rect 79 163 87 171
rect 92 163 100 171
rect 24 64 30 70
rect 13 16 19 22
rect 23 -59 29 -53
rect 67 -66 75 -58
rect 87 -73 95 -65
rect 9 -104 15 -98
<< psubstratepcontact >>
rect 23 326 30 330
rect 44 326 51 330
rect 66 326 73 330
rect 9 109 16 121
rect 37 109 44 121
rect 66 109 73 121
rect 23 -113 30 -109
rect 60 -113 67 -109
rect 81 -113 88 -109
<< nsubstratencontact >>
rect 12 218 19 229
rect 37 218 44 229
rect 75 218 82 229
rect 11 -5 18 6
rect 36 -5 43 6
rect 74 -5 81 6
<< labels >>
rlabel metal1 77 66 92 70 0 S1
rlabel polysilicon 85 83 100 91 0 S0
rlabel metal2 91 0 100 230 0 MUXOUT
rlabel metal2 52 -115 60 -58 0 REGIN
rlabel metal2 91 -65 100 163 0 MUXOUT
rlabel m2contact 79 163 87 171 0 ADDSUB
rlabel m2contact 67 268 75 276 0 DIVIN
rlabel metal1 0 -115 23 -107 0 GND
rlabel metal1 43 -8 74 8 0 Vdd
<< end >>
