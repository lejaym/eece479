magic
tech scmos
timestamp 1427941508
<< pwell >>
rect -21 -23 18 -1
<< nwell >>
rect -21 2 18 33
<< polysilicon >>
rect -12 25 -10 27
rect -2 25 0 27
rect 8 25 10 27
rect -12 2 -10 5
rect -12 -5 -10 -2
rect -2 -5 0 5
rect 8 -5 10 5
rect -12 -17 -10 -15
rect -2 -23 0 -15
rect 8 -23 10 -15
<< ndiffusion >>
rect -14 -15 -12 -5
rect -10 -15 -8 -5
rect -4 -15 -2 -5
rect 0 -15 2 -5
rect 6 -15 8 -5
rect 10 -15 12 -5
<< pdiffusion >>
rect -14 5 -12 25
rect -10 5 -8 25
rect -4 5 -2 25
rect 0 5 2 25
rect 6 5 8 25
rect 10 5 12 25
<< metal1 >>
rect -21 29 -16 33
rect -6 29 18 33
rect -8 25 -4 29
rect -20 5 -18 9
rect -20 2 -16 5
rect 12 2 16 5
rect -21 -2 -16 2
rect -9 -2 16 2
rect -20 -5 -16 -2
rect 2 -5 6 -2
rect -20 -9 -18 -5
rect -8 -19 -4 -15
rect 12 -19 16 -15
rect -21 -23 -16 -19
rect -6 -23 18 -19
<< ntransistor >>
rect -12 -15 -10 -5
rect -2 -15 0 -5
rect 8 -15 10 -5
<< ptransistor >>
rect -12 5 -10 25
rect -2 5 0 25
rect 8 5 10 25
<< polycontact >>
rect -13 -2 -9 2
<< ndcontact >>
rect -18 -15 -14 -5
rect -8 -15 -4 -5
rect 2 -15 6 -5
rect 12 -15 16 -5
<< pdcontact >>
rect -18 5 -14 25
rect -8 5 -4 25
rect 2 5 6 25
rect 12 5 16 25
<< psubstratepcontact >>
rect -16 -23 -6 -19
<< nsubstratencontact >>
rect -16 29 -6 33
<< labels >>
rlabel metal1 -20 -5 -16 5 3 AorB
rlabel polysilicon 8 -5 10 5 1 B
rlabel polysilicon -2 -5 0 5 1 A
rlabel metal1 -6 29 18 33 5 Vdd
rlabel metal1 -6 -23 18 -19 1 Gnd
<< end >>
