magic
tech scmos
timestamp 1427935691
<< pwell >>
rect -20 -23 10 -2
<< nwell >>
rect -20 2 10 32
<< polysilicon >>
rect -11 25 -9 27
rect -1 25 1 27
rect -11 -5 -9 5
rect -1 -5 1 5
rect -11 -23 -9 -15
rect -1 -23 1 -15
<< ndiffusion >>
rect -13 -15 -11 -5
rect -9 -15 -7 -5
rect -3 -15 -1 -5
rect 1 -15 3 -5
<< pdiffusion >>
rect -13 5 -11 25
rect -9 5 -7 25
rect -3 5 -1 25
rect 1 5 3 25
<< metal1 >>
rect -20 29 -10 33
rect 0 29 10 33
rect -17 25 -13 29
rect 3 25 7 29
rect -7 2 -3 5
rect -20 -2 7 2
rect 3 -5 7 -2
rect -17 -19 -13 -15
rect -20 -23 -8 -19
rect -2 -23 10 -19
<< ntransistor >>
rect -11 -15 -9 -5
rect -1 -15 1 -5
<< ptransistor >>
rect -11 5 -9 25
rect -1 5 1 25
<< ndcontact >>
rect -17 -15 -13 -5
rect -7 -15 -3 -5
rect 3 -15 7 -5
<< pdcontact >>
rect -17 5 -13 25
rect -7 5 -3 25
rect 3 5 7 25
<< psubstratepcontact >>
rect -8 -23 -2 -19
<< nsubstratencontact >>
rect -10 29 0 33
<< labels >>
rlabel polysilicon -1 -5 1 5 1 B
rlabel polysilicon -11 -5 -9 5 1 A
rlabel metal1 0 29 10 33 6 Vdd
rlabel metal1 -2 -23 10 -19 1 Gnd
rlabel metal1 -20 -2 -3 2 1 Out
<< end >>
